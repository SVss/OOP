�� sr java.util.ArrayListx����a� I sizexp   w   sr Instruments.Shapes.Circle�����~  xr Instruments.Shapes.Rectangle�M_)�B;�  xr Instruments.Shapes.RectShape�FVv� L 
firstPointt LInstruments/Shapes/Point;L secondPointq ~ xr Instruments.Shapes.Shape_�6�wא L borderColort Ljava/awt/Color;xpsr java.awt.Color���3u F falphaI valueL cst Ljava/awt/color/ColorSpace;[ 	frgbvaluet [F[ fvalueq ~ xp    �   pppsr Instruments.Shapes.Point)�?5��� I xI yxp  �   �sq ~      �sr Instruments.Shapes.PolyLineE�vY���  xr Instruments.Shapes.PolyShape�\�)���y L 
pointsListt Ljava/util/ArrayList;xq ~ q ~ sq ~     w   sq ~   �   �sq ~   �   ?sq ~      �sq ~   r   �sq ~      ysq ~   �   �xsq ~ sq ~ 	    �   pppsq ~      �sq ~      �sq ~ q ~ sq ~   �   �sq ~   �   �sq ~ q ~ sq ~   a   jsq ~   o   �sq ~ q ~ sq ~      bsq ~   #   ~sq ~ q ~ sq ~   �   /sq ~   �   Esr Instruments.Shapes.EllipseJ|�irES�  xq ~ q ~ sq ~   d   Ssq ~   l   gsq ~ +q ~ sq ~   �   sq ~   �   +sq ~ +q ~ sq ~      �sq ~      �sq ~ +q ~ sq ~      Osq ~      asq ~ +q ~ sq ~   �   �sq ~   �   �x